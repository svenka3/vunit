-- This Source Code Form is subject to the terms of the Mozilla Public
-- License, v. 2.0. If a copy of the MPL was not distributed with this file,
-- You can obtain one at http://mozilla.org/MPL/2.0/.
--
-- Copyright (c) 2016, Lars Asplund lars.anders.asplund@gmail.com

package array_assert_pkg is
  procedure array_assert (condition : boolean; msg : string := "");
end package;

package body array_assert_pkg is
  procedure array_assert (condition : boolean; msg : string := "") is
  begin
    assert condition report msg;
  end;
end package body array_assert_pkg;
